`include "quadra.vh"

module lut
(
    input  x1_t  x1,
    output a_t   a,
    output b_t   b,
    output c_t   c
);
    // Read coefficients:
    always_comb
    unique casez (x1)
        7'b0000000 :  a = 24'ha57d87;
        7'b0000001 :  a = 24'ha85ccc;
        7'b0000010 :  a = 24'hab51fb;
        7'b0000011 :  a = 24'hae5c54;
        7'b0000100 :  a = 24'hb17b15;
        7'b0000101 :  a = 24'hb4ad78;
        7'b0000110 :  a = 24'hb7f2ae;
        7'b0000111 :  a = 24'hbb49e8;
        7'b0001000 :  a = 24'hbeb24e;
        7'b0001001 :  a = 24'hc22b09;
        7'b0001010 :  a = 24'hc5b337;
        7'b0001011 :  a = 24'hc949f9;
        7'b0001100 :  a = 24'hccee68;
        7'b0001101 :  a = 24'hd09f9b;
        7'b0001110 :  a = 24'hd45ca6;
        7'b0001111 :  a = 24'hd82499;
        7'b0010000 :  a = 24'hdbf683;
        7'b0010001 :  a = 24'hdfd170;
        7'b0010010 :  a = 24'he3b468;
        7'b0010011 :  a = 24'he79e72;
        7'b0010100 :  a = 24'heb8e95;
        7'b0010101 :  a = 24'hef83d4;
        7'b0010110 :  a = 24'hf37d32;
        7'b0010111 :  a = 24'hf779b1;
        7'b0011000 :  a = 24'hfb7851;
        7'b0011001 :  a = 24'hff7813;
        7'b0011010 :  a = 24'h0377f6;
        7'b0011011 :  a = 24'h0776fc;
        7'b0011100 :  a = 24'h0b7425;
        7'b0011101 :  a = 24'h0f6e70;
        7'b0011110 :  a = 24'h1364e0;
        7'b0011111 :  a = 24'h175677;
        7'b0100000 :  a = 24'h1b4238;
        7'b0100001 :  a = 24'h1f2729;
        7'b0100010 :  a = 24'h230450;
        7'b0100011 :  a = 24'h26d8b6;
        7'b0100100 :  a = 24'h2aa367;
        7'b0100101 :  a = 24'h2e636e;
        7'b0100110 :  a = 24'h3217de;
        7'b0100111 :  a = 24'h35bfc7;
        7'b0101000 :  a = 24'h395a41;
        7'b0101001 :  a = 24'h3ce664;
        7'b0101010 :  a = 24'h40634e;
        7'b0101011 :  a = 24'h43d020;
        7'b0101100 :  a = 24'h472bfe;
        7'b0101101 :  a = 24'h4a7611;
        7'b0101110 :  a = 24'h4dad88;
        7'b0101111 :  a = 24'h50d193;
        7'b0110000 :  a = 24'h53e16b;
        7'b0110001 :  a = 24'h56dc4a;
        7'b0110010 :  a = 24'h59c173;
        7'b0110011 :  a = 24'h5c902b;
        7'b0110100 :  a = 24'h5f47c1;
        7'b0110101 :  a = 24'h61e785;
        7'b0110110 :  a = 24'h646ecf;
        7'b0110111 :  a = 24'h66dcff;
        7'b0111000 :  a = 24'h693177;
        7'b0111001 :  a = 24'h6b6ba4;
        7'b0111010 :  a = 24'h6d8af6;
        7'b0111011 :  a = 24'h6f8ee7;
        7'b0111100 :  a = 24'h7176f4;
        7'b0111101 :  a = 24'h7342a4;
        7'b0111110 :  a = 24'h74f184;
        7'b0111111 :  a = 24'h768328;
        7'b1000000 :  a = 24'h77f72c;
        7'b1000001 :  a = 24'h794d33;
        7'b1000010 :  a = 24'h7a84e7;
        7'b1000011 :  a = 24'h7b9dfa;
        7'b1000100 :  a = 24'h7c9827;
        7'b1000101 :  a = 24'h7d732e;
        7'b1000110 :  a = 24'h7e2ed9;
        7'b1000111 :  a = 24'h7ecafa;
        7'b1001000 :  a = 24'h7f4768;
        7'b1001001 :  a = 24'h7fa405;
        7'b1001010 :  a = 24'h7fe0b9;
        7'b1001011 :  a = 24'h7ffd76;
        7'b1001100 :  a = 24'h7ffa34;
        7'b1001101 :  a = 24'h7fd6f5;
        7'b1001110 :  a = 24'h7f93c0;
        7'b1001111 :  a = 24'h7f30a7;
        7'b1010000 :  a = 24'h7eadc3;
        7'b1010001 :  a = 24'h7e0b33;
        7'b1010010 :  a = 24'h7d4922;
        7'b1010011 :  a = 24'h7c67bf;
        7'b1010100 :  a = 24'h7b6743;
        7'b1010101 :  a = 24'h7a47ed;
        7'b1010110 :  a = 24'h790a07;
        7'b1010111 :  a = 24'h77adde;
        7'b1011000 :  a = 24'h7633ca;
        7'b1011001 :  a = 24'h749c2a;
        7'b1011010 :  a = 24'h72e764;
        7'b1011011 :  a = 24'h7115e5;
        7'b1011100 :  a = 24'h6f2820;
        7'b1011101 :  a = 24'h6d1e92;
        7'b1011110 :  a = 24'h6af9bd;
        7'b1011111 :  a = 24'h68ba2b;
        7'b1100000 :  a = 24'h66606a;
        7'b1100001 :  a = 24'h63ed11;
        7'b1100010 :  a = 24'h6160be;
        7'b1100011 :  a = 24'h5ebc13;
        7'b1100100 :  a = 24'h5bffba;
        7'b1100101 :  a = 24'h592c61;
        7'b1100110 :  a = 24'h5642be;
        7'b1100111 :  a = 24'h53438a;
        7'b1101000 :  a = 24'h502f86;
        7'b1101001 :  a = 24'h4d0777;
        7'b1101010 :  a = 24'h49cc25;
        7'b1101011 :  a = 24'h467e62;
        7'b1101100 :  a = 24'h431eff;
        7'b1101101 :  a = 24'h3faed4;
        7'b1101110 :  a = 24'h3c2ebf;
        7'b1101111 :  a = 24'h389f9e;
        7'b1110000 :  a = 24'h350255;
        7'b1110001 :  a = 24'h3157cc;
        7'b1110010 :  a = 24'h2da0ed;
        7'b1110011 :  a = 24'h29dea7;
        7'b1110100 :  a = 24'h2611e8;
        7'b1110101 :  a = 24'h223ba6;
        7'b1110110 :  a = 24'h1e5cd5;
        7'b1110111 :  a = 24'h1a766d;
        7'b1111000 :  a = 24'h168967;
        7'b1111001 :  a = 24'h1296bf;
        7'b1111010 :  a = 24'h0e9f72;
        7'b1111011 :  a = 24'h0aa47c;
        7'b1111100 :  a = 24'h06a6de;
        7'b1111101 :  a = 24'h02a796;
        7'b1111110 :  a = 24'hfea7a5;
        7'b1111111 :  a = 24'hfaa809;
        default    :  a = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  b = 19'h16a0c;
        7'b0000001 :  b = 19'h1752f;
        7'b0000010 :  b = 19'h17ff4;
        7'b0000011 :  b = 19'h18a59;
        7'b0000100 :  b = 19'h1945c;
        7'b0000101 :  b = 19'h19dfa;
        7'b0000110 :  b = 19'h1a730;
        7'b0000111 :  b = 19'h1affd;
        7'b0001000 :  b = 19'h1b85d;
        7'b0001001 :  b = 19'h1c04f;
        7'b0001010 :  b = 19'h1c7d2;
        7'b0001011 :  b = 19'h1cee2;
        7'b0001100 :  b = 19'h1d57f;
        7'b0001101 :  b = 19'h1dba6;
        7'b0001110 :  b = 19'h1e156;
        7'b0001111 :  b = 19'h1e68e;
        7'b0010000 :  b = 19'h1eb4d;
        7'b0010001 :  b = 19'h1ef91;
        7'b0010010 :  b = 19'h1f358;
        7'b0010011 :  b = 19'h1f6a3;
        7'b0010100 :  b = 19'h1f970;
        7'b0010101 :  b = 19'h1fbbf;
        7'b0010110 :  b = 19'h1fd8f;
        7'b0010111 :  b = 19'h1fee0;
        7'b0011000 :  b = 19'h1ffb1;
        7'b0011001 :  b = 19'h20002;
        7'b0011010 :  b = 19'h1ffd3;
        7'b0011011 :  b = 19'h1ff24;
        7'b0011100 :  b = 19'h1fdf5;
        7'b0011101 :  b = 19'h1fc47;
        7'b0011110 :  b = 19'h1fa1a;
        7'b0011111 :  b = 19'h1f76e;
        7'b0100000 :  b = 19'h1f444;
        7'b0100001 :  b = 19'h1f09e;
        7'b0100010 :  b = 19'h1ec7b;
        7'b0100011 :  b = 19'h1e7dd;
        7'b0100100 :  b = 19'h1e2c5;
        7'b0100101 :  b = 19'h1dd34;
        7'b0100110 :  b = 19'h1d72c;
        7'b0100111 :  b = 19'h1d0af;
        7'b0101000 :  b = 19'h1c9bd;
        7'b0101001 :  b = 19'h1c259;
        7'b0101010 :  b = 19'h1ba84;
        7'b0101011 :  b = 19'h1b240;
        7'b0101100 :  b = 19'h1a990;
        7'b0101101 :  b = 19'h1a076;
        7'b0101110 :  b = 19'h196f4;
        7'b0101111 :  b = 19'h18d0b;
        7'b0110000 :  b = 19'h182c0;
        7'b0110001 :  b = 19'h17814;
        7'b0110010 :  b = 19'h16d0a;
        7'b0110011 :  b = 19'h161a4;
        7'b0110100 :  b = 19'h155e6;
        7'b0110101 :  b = 19'h149d3;
        7'b0110110 :  b = 19'h13d6d;
        7'b0110111 :  b = 19'h130b8;
        7'b0111000 :  b = 19'h123b7;
        7'b0111001 :  b = 19'h1166d;
        7'b0111010 :  b = 19'h108dd;
        7'b0111011 :  b = 19'h0fb0b;
        7'b0111100 :  b = 19'h0ecfa;
        7'b0111101 :  b = 19'h0deae;
        7'b0111110 :  b = 19'h0d02b;
        7'b0111111 :  b = 19'h0c173;
        7'b1000000 :  b = 19'h0b28b;
        7'b1000001 :  b = 19'h0a376;
        7'b1000010 :  b = 19'h09439;
        7'b1000011 :  b = 19'h084d6;
        7'b1000100 :  b = 19'h07552;
        7'b1000101 :  b = 19'h065b1;
        7'b1000110 :  b = 19'h055f7;
        7'b1000111 :  b = 19'h04627;
        7'b1001000 :  b = 19'h03645;
        7'b1001001 :  b = 19'h02656;
        7'b1001010 :  b = 19'h0165d;
        7'b1001011 :  b = 19'h0065f;
        7'b1001100 :  b = 19'h7f65f;
        7'b1001101 :  b = 19'h7e662;
        7'b1001110 :  b = 19'h7d66b;
        7'b1001111 :  b = 19'h7c67e;
        7'b1010000 :  b = 19'h7b6a0;
        7'b1010001 :  b = 19'h7a6d4;
        7'b1010010 :  b = 19'h7971e;
        7'b1010011 :  b = 19'h78783;
        7'b1010100 :  b = 19'h77805;
        7'b1010101 :  b = 19'h768aa;
        7'b1010110 :  b = 19'h75974;
        7'b1010111 :  b = 19'h74a68;
        7'b1011000 :  b = 19'h73b8a;
        7'b1011001 :  b = 19'h72cdd;
        7'b1011010 :  b = 19'h71e64;
        7'b1011011 :  b = 19'h71024;
        7'b1011100 :  b = 19'h7021f;
        7'b1011101 :  b = 19'h6f45b;
        7'b1011110 :  b = 19'h6e6d9;
        7'b1011111 :  b = 19'h6d99d;
        7'b1100000 :  b = 19'h6ccab;
        7'b1100001 :  b = 19'h6c006;
        7'b1100010 :  b = 19'h6b3b1;
        7'b1100011 :  b = 19'h6a7af;
        7'b1100100 :  b = 19'h69c03;
        7'b1100101 :  b = 19'h690b0;
        7'b1100110 :  b = 19'h685b8;
        7'b1100111 :  b = 19'h67b20;
        7'b1101000 :  b = 19'h670e8;
        7'b1101001 :  b = 19'h66714;
        7'b1101010 :  b = 19'h65da7;
        7'b1101011 :  b = 19'h654a2;
        7'b1101100 :  b = 19'h64c08;
        7'b1101101 :  b = 19'h643db;
        7'b1101110 :  b = 19'h63c1d;
        7'b1101111 :  b = 19'h634d0;
        7'b1110000 :  b = 19'h62df5;
        7'b1110001 :  b = 19'h62790;
        7'b1110010 :  b = 19'h621a0;
        7'b1110011 :  b = 19'h61c28;
        7'b1110100 :  b = 19'h61729;
        7'b1110101 :  b = 19'h612a4;
        7'b1110110 :  b = 19'h60e9a;
        7'b1110111 :  b = 19'h60b0d;
        7'b1111000 :  b = 19'h607fd;
        7'b1111001 :  b = 19'h6056b;
        7'b1111010 :  b = 19'h60357;
        7'b1111011 :  b = 19'h601c3;
        7'b1111100 :  b = 19'h600ae;
        7'b1111101 :  b = 19'h60019;
        7'b1111110 :  b = 19'h60004;
        7'b1111111 :  b = 19'h6006f;
        default    :  b = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  c = 13'h0b39;
        7'b0000001 :  c = 13'h0add;
        7'b0000010 :  c = 13'h0a7d;
        7'b0000011 :  c = 13'h0a1b;
        7'b0000100 :  c = 13'h09b7;
        7'b0000101 :  c = 13'h0950;
        7'b0000110 :  c = 13'h08e7;
        7'b0000111 :  c = 13'h087b;
        7'b0001000 :  c = 13'h080e;
        7'b0001001 :  c = 13'h079e;
        7'b0001010 :  c = 13'h072d;
        7'b0001011 :  c = 13'h06ba;
        7'b0001100 :  c = 13'h0645;
        7'b0001101 :  c = 13'h05ce;
        7'b0001110 :  c = 13'h0556;
        7'b0001111 :  c = 13'h04dd;
        7'b0010000 :  c = 13'h0462;
        7'b0010001 :  c = 13'h03e7;
        7'b0010010 :  c = 13'h036a;
        7'b0010011 :  c = 13'h02ed;
        7'b0010100 :  c = 13'h026e;
        7'b0010101 :  c = 13'h01f0;
        7'b0010110 :  c = 13'h0170;
        7'b0010111 :  c = 13'h00f1;
        7'b0011000 :  c = 13'h0071;
        7'b0011001 :  c = 13'h1ff1;
        7'b0011010 :  c = 13'h1f71;
        7'b0011011 :  c = 13'h1ef1;
        7'b0011100 :  c = 13'h1e72;
        7'b0011101 :  c = 13'h1df3;
        7'b0011110 :  c = 13'h1d74;
        7'b0011111 :  c = 13'h1cf6;
        7'b0100000 :  c = 13'h1c79;
        7'b0100001 :  c = 13'h1bfc;
        7'b0100010 :  c = 13'h1b81;
        7'b0100011 :  c = 13'h1b07;
        7'b0100100 :  c = 13'h1a8e;
        7'b0100101 :  c = 13'h1a16;
        7'b0100110 :  c = 13'h19a0;
        7'b0100111 :  c = 13'h192b;
        7'b0101000 :  c = 13'h18b8;
        7'b0101001 :  c = 13'h1847;
        7'b0101010 :  c = 13'h17d8;
        7'b0101011 :  c = 13'h176b;
        7'b0101100 :  c = 13'h1700;
        7'b0101101 :  c = 13'h1698;
        7'b0101110 :  c = 13'h1631;
        7'b0101111 :  c = 13'h15cd;
        7'b0110000 :  c = 13'h156c;
        7'b0110001 :  c = 13'h150d;
        7'b0110010 :  c = 13'h14b1;
        7'b0110011 :  c = 13'h1458;
        7'b0110100 :  c = 13'h1402;
        7'b0110101 :  c = 13'h13af;
        7'b0110110 :  c = 13'h135f;
        7'b0110111 :  c = 13'h1312;
        7'b0111000 :  c = 13'h12c8;
        7'b0111001 :  c = 13'h1282;
        7'b0111010 :  c = 13'h123e;
        7'b0111011 :  c = 13'h11ff;
        7'b0111100 :  c = 13'h11c3;
        7'b0111101 :  c = 13'h118a;
        7'b0111110 :  c = 13'h1155;
        7'b0111111 :  c = 13'h1124;
        7'b1000000 :  c = 13'h10f6;
        7'b1000001 :  c = 13'h10cd;
        7'b1000010 :  c = 13'h10a7;
        7'b1000011 :  c = 13'h1084;
        7'b1000100 :  c = 13'h1066;
        7'b1000101 :  c = 13'h104c;
        7'b1000110 :  c = 13'h1035;
        7'b1000111 :  c = 13'h1023;
        7'b1001000 :  c = 13'h1014;
        7'b1001001 :  c = 13'h1009;
        7'b1001010 :  c = 13'h1003;
        7'b1001011 :  c = 13'h1000;
        7'b1001100 :  c = 13'h1002;
        7'b1001101 :  c = 13'h1007;
        7'b1001110 :  c = 13'h1011;
        7'b1001111 :  c = 13'h101e;
        7'b1010000 :  c = 13'h102f;
        7'b1010001 :  c = 13'h1045;
        7'b1010010 :  c = 13'h105e;
        7'b1010011 :  c = 13'h107b;
        7'b1010100 :  c = 13'h109c;
        7'b1010101 :  c = 13'h10c1;
        7'b1010110 :  c = 13'h10ea;
        7'b1010111 :  c = 13'h1116;
        7'b1011000 :  c = 13'h1146;
        7'b1011001 :  c = 13'h117a;
        7'b1011010 :  c = 13'h11b2;
        7'b1011011 :  c = 13'h11ed;
        7'b1011100 :  c = 13'h122b;
        7'b1011101 :  c = 13'h126d;
        7'b1011110 :  c = 13'h12b3;
        7'b1011111 :  c = 13'h12fb;
        7'b1100000 :  c = 13'h1348;
        7'b1100001 :  c = 13'h1397;
        7'b1100010 :  c = 13'h13e9;
        7'b1100011 :  c = 13'h143e;
        7'b1100100 :  c = 13'h1497;
        7'b1100101 :  c = 13'h14f2;
        7'b1100110 :  c = 13'h1550;
        7'b1100111 :  c = 13'h15b0;
        7'b1101000 :  c = 13'h1613;
        7'b1101001 :  c = 13'h1679;
        7'b1101010 :  c = 13'h16e1;
        7'b1101011 :  c = 13'h174b;
        7'b1101100 :  c = 13'h17b8;
        7'b1101101 :  c = 13'h1826;
        7'b1101110 :  c = 13'h1897;
        7'b1101111 :  c = 13'h1909;
        7'b1110000 :  c = 13'h197d;
        7'b1110001 :  c = 13'h19f3;
        7'b1110010 :  c = 13'h1a6a;
        7'b1110011 :  c = 13'h1ae3;
        7'b1110100 :  c = 13'h1b5d;
        7'b1110101 :  c = 13'h1bd8;
        7'b1110110 :  c = 13'h1c54;
        7'b1110111 :  c = 13'h1cd1;
        7'b1111000 :  c = 13'h1d4f;
        7'b1111001 :  c = 13'h1dcd;
        7'b1111010 :  c = 13'h1e4c;
        7'b1111011 :  c = 13'h1ecc;
        7'b1111100 :  c = 13'h1f4b;
        7'b1111101 :  c = 13'h1fcb;
        7'b1111110 :  c = 13'h004b;
        7'b1111111 :  c = 13'h00cb;
        default    :  c = 'x;
    endcase

endmodule
