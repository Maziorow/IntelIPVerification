`include "quadra.vh"

module lut
(
    input  x1_t  x1,
    output a_t   a,
    output b_t   b,
    output c_t   c
);
    // Read coefficients:
    always_comb
    unique casez (x1)
        7'b0000000 :  a = 32'hf4afb0cd;
        7'b0000001 :  a = 32'hf50b9983;
        7'b0000010 :  a = 32'hf56a3f45;
        7'b0000011 :  a = 32'hf5cb8a69;
        7'b0000100 :  a = 32'hf62f629c;
        7'b0000101 :  a = 32'hf695aeea;
        7'b0000110 :  a = 32'hf6fe55bf;
        7'b0000111 :  a = 32'hf7693cf3;
        7'b0001000 :  a = 32'hf7d649cc;
        7'b0001001 :  a = 32'hf8456108;
        7'b0001010 :  a = 32'hf8b666e2;
        7'b0001011 :  a = 32'hf9293f18;
        7'b0001100 :  a = 32'hf99dccf5;
        7'b0001101 :  a = 32'hfa13f356;
        7'b0001110 :  a = 32'hfa8b94b3;
        7'b0001111 :  a = 32'hfb049323;
        7'b0010000 :  a = 32'hfb7ed068;
        7'b0010001 :  a = 32'hfbfa2df2;
        7'b0010010 :  a = 32'hfc768cec;
        7'b0010011 :  a = 32'hfcf3ce3e;
        7'b0010100 :  a = 32'hfd71d298;
        7'b0010101 :  a = 32'hfdf07a7a;
        7'b0010110 :  a = 32'hfe6fa63b;
        7'b0010111 :  a = 32'hfeef3610;
        7'b0011000 :  a = 32'hff6f0a16;
        7'b0011001 :  a = 32'hffef0259;
        7'b0011010 :  a = 32'h006efedb;
        7'b0011011 :  a = 32'h00eedf9e;
        7'b0011100 :  a = 32'h016e84ab;
        7'b0011101 :  a = 32'h01edce18;
        7'b0011110 :  a = 32'h026c9c14;
        7'b0011111 :  a = 32'h02eaceed;
        7'b0100000 :  a = 32'h03684715;
        7'b0100001 :  a = 32'h03e4e531;
        7'b0100010 :  a = 32'h04608a18;
        7'b0100011 :  a = 32'h04db16e2;
        7'b0100100 :  a = 32'h05546cee;
        7'b0100101 :  a = 32'h05cc6de5;
        7'b0100110 :  a = 32'h0642fbc8;
        7'b0100111 :  a = 32'h06b7f8f5;
        7'b0101000 :  a = 32'h072b482d;
        7'b0101001 :  a = 32'h079ccc9c;
        7'b0101010 :  a = 32'h080c69e2;
        7'b0101011 :  a = 32'h087a0419;
        7'b0101100 :  a = 32'h08e57fd9;
        7'b0101101 :  a = 32'h094ec246;
        7'b0101110 :  a = 32'h09b5b10e;
        7'b0101111 :  a = 32'h0a1a3277;
        7'b0110000 :  a = 32'h0a7c2d61;
        7'b0110001 :  a = 32'h0adb894e;
        7'b0110010 :  a = 32'h0b382e66;
        7'b0110011 :  a = 32'h0b920582;
        7'b0110100 :  a = 32'h0be8f82c;
        7'b0110101 :  a = 32'h0c3cf0a8;
        7'b0110110 :  a = 32'h0c8dd9f8;
        7'b0110111 :  a = 32'h0cdb9fe3;
        7'b0111000 :  a = 32'h0d262ef6;
        7'b0111001 :  a = 32'h0d6d7490;
        7'b0111010 :  a = 32'h0db15ede;
        7'b0111011 :  a = 32'h0df1dce6;
        7'b0111100 :  a = 32'h0e2ede8a;
        7'b0111101 :  a = 32'h0e685489;
        7'b0111110 :  a = 32'h0e9e3087;
        7'b0111111 :  a = 32'h0ed0650b;
        7'b1000000 :  a = 32'h0efee58b;
        7'b1000001 :  a = 32'h0f29a664;
        7'b1000010 :  a = 32'h0f509ce9;
        7'b1000011 :  a = 32'h0f73bf5a;
        7'b1000100 :  a = 32'h0f9304f1;
        7'b1000101 :  a = 32'h0fae65db;
        7'b1000110 :  a = 32'h0fc5db40;
        7'b1000111 :  a = 32'h0fd95f44;
        7'b1001000 :  a = 32'h0fe8ed04;
        7'b1001001 :  a = 32'h0ff4809f;
        7'b1001010 :  a = 32'h0ffc172f;
        7'b1001011 :  a = 32'h0fffaecf;
        7'b1001100 :  a = 32'h0fff4698;
        7'b1001101 :  a = 32'h0ffadea4;
        7'b1001110 :  a = 32'h0ff2780f;
        7'b1001111 :  a = 32'h0fe614f0;
        7'b1010000 :  a = 32'h0fd5b862;
        7'b1010001 :  a = 32'h0fc1667b;
        7'b1010010 :  a = 32'h0fa9244f;
        7'b1010011 :  a = 32'h0f8cf7ef;
        7'b1010100 :  a = 32'h0f6ce865;
        7'b1010101 :  a = 32'h0f48fdb6;
        7'b1010110 :  a = 32'h0f2140dc;
        7'b1010111 :  a = 32'h0ef5bbc6;
        7'b1011000 :  a = 32'h0ec67955;
        7'b1011001 :  a = 32'h0e938559;
        7'b1011010 :  a = 32'h0e5cec90;
        7'b1011011 :  a = 32'h0e22bc9e;
        7'b1011100 :  a = 32'h0de50410;
        7'b1011101 :  a = 32'h0da3d254;
        7'b1011110 :  a = 32'h0d5f37b5;
        7'b1011111 :  a = 32'h0d17455a;
        7'b1100000 :  a = 32'h0ccc0d40;
        7'b1100001 :  a = 32'h0c7da233;
        7'b1100010 :  a = 32'h0c2c17ce;
        7'b1100011 :  a = 32'h0bd78273;
        7'b1100100 :  a = 32'h0b7ff748;
        7'b1100101 :  a = 32'h0b258c2e;
        7'b1100110 :  a = 32'h0ac857c0;
        7'b1100111 :  a = 32'h0a68714a;
        7'b1101000 :  a = 32'h0a05f0c6;
        7'b1101001 :  a = 32'h09a0eed3;
        7'b1101010 :  a = 32'h093984b1;
        7'b1101011 :  a = 32'h08cfcc3a;
        7'b1101100 :  a = 32'h0863dfdc;
        7'b1101101 :  a = 32'h07f5da92;
        7'b1101110 :  a = 32'h0785d7db;
        7'b1101111 :  a = 32'h0713f3b8;
        7'b1110000 :  a = 32'h06a04aa2;
        7'b1110001 :  a = 32'h062af982;
        7'b1110010 :  a = 32'h05b41dac;
        7'b1110011 :  a = 32'h053bd4d6;
        7'b1110100 :  a = 32'h04c23d11;
        7'b1110101 :  a = 32'h044774c4;
        7'b1110110 :  a = 32'h03cb9a9f;
        7'b1110111 :  a = 32'h034ecd99;
        7'b1111000 :  a = 32'h02d12ce4;
        7'b1111001 :  a = 32'h0252d7e7;
        7'b1111010 :  a = 32'h01d3ee38;
        7'b1111011 :  a = 32'h01548f8f;
        7'b1111100 :  a = 32'h00d4dbc4;
        7'b1111101 :  a = 32'h0054f2c3;
        7'b1111110 :  a = 32'hffd4f487;
        7'b1111111 :  a = 32'hff55010c;
        default    :  a = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  b = 32'h16a09e66;
        7'b0000001 :  b = 32'h1752c7ca;
        7'b0000010 :  b = 32'h17ff1c9b;
        7'b0000011 :  b = 32'h18a571c5;
        7'b0000100 :  b = 32'h19459db3;
        7'b0000101 :  b = 32'h19df785b;
        7'b0000110 :  b = 32'h1a72db48;
        7'b0000111 :  b = 32'h1affa1a1;
        7'b0001000 :  b = 32'h1b85a836;
        7'b0001001 :  b = 32'h1c04cd86;
        7'b0001010 :  b = 32'h1c7cf1c7;
        7'b0001011 :  b = 32'h1cedf6f2;
        7'b0001100 :  b = 32'h1d57c0c6;
        7'b0001101 :  b = 32'h1dba34d1;
        7'b0001110 :  b = 32'h1e153a76;
        7'b0001111 :  b = 32'h1e68baf4;
        7'b0010000 :  b = 32'h1eb4a16d;
        7'b0010001 :  b = 32'h1ef8dae6;
        7'b0010010 :  b = 32'h1f355652;
        7'b0010011 :  b = 32'h1f6a0491;
        7'b0010100 :  b = 32'h1f96d87a;
        7'b0010101 :  b = 32'h1fbbc6d6;
        7'b0010110 :  b = 32'h1fd8c66b;
        7'b0010111 :  b = 32'h1fedcff9;
        7'b0011000 :  b = 32'h1ffade3d;
        7'b0011001 :  b = 32'h1fffedf5;
        7'b0011010 :  b = 32'h1ffcfddc;
        7'b0011011 :  b = 32'h1ff20eae;
        7'b0011100 :  b = 32'h1fdf2326;
        7'b0011101 :  b = 32'h1fc44001;
        7'b0011110 :  b = 32'h1fa16bf6;
        7'b0011111 :  b = 32'h1f76afba;
        7'b0100000 :  b = 32'h1f4415fc;
        7'b0100001 :  b = 32'h1f09ab62;
        7'b0100010 :  b = 32'h1ec77e87;
        7'b0100011 :  b = 32'h1e7d9ff5;
        7'b0100100 :  b = 32'h1e2c2224;
        7'b0100101 :  b = 32'h1dd31972;
        7'b0100110 :  b = 32'h1d729c22;
        7'b0100111 :  b = 32'h1d0ac253;
        7'b0101000 :  b = 32'h1c9ba5f9;
        7'b0101001 :  b = 32'h1c2562dc;
        7'b0101010 :  b = 32'h1ba8168c;
        7'b0101011 :  b = 32'h1b23e05b;
        7'b0101100 :  b = 32'h1a98e156;
        7'b0101101 :  b = 32'h1a073c3c;
        7'b0101110 :  b = 32'h196f1576;
        7'b0101111 :  b = 32'h18d0930c;
        7'b0110000 :  b = 32'h182bdc9f;
        7'b0110001 :  b = 32'h17811b5b;
        7'b0110010 :  b = 32'h16d079ef;
        7'b0110011 :  b = 32'h161a2484;
        7'b0110100 :  b = 32'h155e48ac;
        7'b0110101 :  b = 32'h149d155f;
        7'b0110110 :  b = 32'h13d6bae8;
        7'b0110111 :  b = 32'h130b6add;
        7'b0111000 :  b = 32'h123b5811;
        7'b0111001 :  b = 32'h1166b686;
        7'b0111010 :  b = 32'h108dbb66;
        7'b0111011 :  b = 32'h0fb09cec;
        7'b0111100 :  b = 32'h0ecf9260;
        7'b0111101 :  b = 32'h0dead404;
        7'b0111110 :  b = 32'h0d029b05;
        7'b0111111 :  b = 32'h0c172170;
        7'b1000000 :  b = 32'h0b28a224;
        7'b1000001 :  b = 32'h0a3758bd;
        7'b1000010 :  b = 32'h0943818e;
        7'b1000011 :  b = 32'h084d598b;
        7'b1000100 :  b = 32'h07551e3d;
        7'b1000101 :  b = 32'h065b0db1;
        7'b1000110 :  b = 32'h055f666a;
        7'b1000111 :  b = 32'h04626751;
        7'b1001000 :  b = 32'h03644fa3;
        7'b1001001 :  b = 32'h02655ee6;
        7'b1001010 :  b = 32'h0165d4d5;
        7'b1001011 :  b = 32'h0065f150;
        7'b1001100 :  b = 32'hff65f450;
        7'b1001101 :  b = 32'hfe661dd1;
        7'b1001110 :  b = 32'hfd66adca;
        7'b1001111 :  b = 32'hfc67e413;
        7'b1010000 :  b = 32'hfb6a005e;
        7'b1010001 :  b = 32'hfa6d4223;
        7'b1010010 :  b = 32'hf971e890;
        7'b1010011 :  b = 32'hf878327b;
        7'b1010100 :  b = 32'hf7805e4e;
        7'b1010101 :  b = 32'hf68aa9ff;
        7'b1010110 :  b = 32'hf59752f8;
        7'b1010111 :  b = 32'hf4a6960f;
        7'b1011000 :  b = 32'hf3b8af72;
        7'b1011001 :  b = 32'hf2cdda98;
        7'b1011010 :  b = 32'hf1e65236;
        7'b1011011 :  b = 32'hf102502c;
        7'b1011100 :  b = 32'hf0220d7b;
        7'b1011101 :  b = 32'hef45c231;
        7'b1011110 :  b = 32'hee6da560;
        7'b1011111 :  b = 32'hed99ed0e;
        7'b1100000 :  b = 32'heccace28;
        7'b1100001 :  b = 32'hec007c76;
        7'b1100010 :  b = 32'heb3b2a89;
        7'b1100011 :  b = 32'hea7b09b7;
        7'b1100100 :  b = 32'he9c04a05;
        7'b1100101 :  b = 32'he90b1a23;
        7'b1100110 :  b = 32'he85ba75c;
        7'b1100111 :  b = 32'he7b21d8b;
        7'b1101000 :  b = 32'he70ea713;
        7'b1101001 :  b = 32'he6716cd0;
        7'b1101010 :  b = 32'he5da960f;
        7'b1101011 :  b = 32'he54a4886;
        7'b1101100 :  b = 32'he4c0a847;
        7'b1101101 :  b = 32'he43dd7ba;
        7'b1101110 :  b = 32'he3c1f792;
        7'b1101111 :  b = 32'he34d26c6;
        7'b1110000 :  b = 32'he2df828b;
        7'b1110001 :  b = 32'he2792648;
        7'b1110010 :  b = 32'he21a2b94;
        7'b1110011 :  b = 32'he1c2aa2d;
        7'b1110100 :  b = 32'he172b7f3;
        7'b1110101 :  b = 32'he12a68e3;
        7'b1110110 :  b = 32'he0e9cf0f;
        7'b1110111 :  b = 32'he0b0fa9f;
        7'b1111000 :  b = 32'he07ff9c5;
        7'b1111001 :  b = 32'he056d8c4;
        7'b1111010 :  b = 32'he035a1e2;
        7'b1111011 :  b = 32'he01c5d6d;
        7'b1111100 :  b = 32'he00b11b6;
        7'b1111101 :  b = 32'he001c310;
        7'b1111110 :  b = 32'he00073cf;
        7'b1111111 :  b = 32'he0072446;
        default    :  b = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  c = 32'h16a09e66;
        7'b0000001 :  c = 32'h15e8ccf9;
        7'b0000010 :  c = 32'h152b8176;
        7'b0000011 :  c = 32'h1468eb2f;
        7'b0000100 :  c = 32'h13a13ac8;
        7'b0000101 :  c = 32'h12d4a22d;
        7'b0000110 :  c = 32'h12035482;
        7'b0000111 :  c = 32'h112d861a;
        7'b0001000 :  c = 32'h10536c67;
        7'b0001001 :  c = 32'h0f753def;
        7'b0001010 :  c = 32'h0e93323c;
        7'b0001011 :  c = 32'h0dad81d1;
        7'b0001100 :  c = 32'h0cc46616;
        7'b0001101 :  c = 32'h0bd81954;
        7'b0001110 :  c = 32'h0ae8d69b;
        7'b0001111 :  c = 32'h09f6d9ba;
        7'b0010000 :  c = 32'h09025f31;
        7'b0010001 :  c = 32'h080ba41c;
        7'b0010010 :  c = 32'h0712e628;
        7'b0010011 :  c = 32'h06186384;
        7'b0010100 :  c = 32'h051c5ad0;
        7'b0010101 :  c = 32'h041f0b0c;
        7'b0010110 :  c = 32'h0320b38a;
        7'b0010111 :  c = 32'h022193e0;
        7'b0011000 :  c = 32'h0121ebd4;
        7'b0011001 :  c = 32'h0021fb4e;
        7'b0011010 :  c = 32'hff220249;
        7'b0011011 :  c = 32'hfe2240c3;
        7'b0011100 :  c = 32'hfd22f6aa;
        7'b0011101 :  c = 32'hfc2463d0;
        7'b0011110 :  c = 32'hfb26c7d8;
        7'b0011111 :  c = 32'hfa2a6227;
        7'b0100000 :  c = 32'hf92f71d5;
        7'b0100001 :  c = 32'hf836359f;
        7'b0100010 :  c = 32'hf73eebd0;
        7'b0100011 :  c = 32'hf649d23b;
        7'b0100100 :  c = 32'hf5572624;
        7'b0100101 :  c = 32'hf4672436;
        7'b0100110 :  c = 32'hf37a086f;
        7'b0100111 :  c = 32'hf2900e15;
        7'b0101000 :  c = 32'hf1a96fa6;
        7'b0101001 :  c = 32'hf0c666c8;
        7'b0101010 :  c = 32'hefe72c3c;
        7'b0101011 :  c = 32'hef0bf7cf;
        7'b0101100 :  c = 32'hee35004e;
        7'b0101101 :  c = 32'hed627b75;
        7'b0101110 :  c = 32'hec949de4;
        7'b0101111 :  c = 32'hebcb9b12;
        7'b0110000 :  c = 32'heb07a53e;
        7'b0110001 :  c = 32'hea48ed65;
        7'b0110010 :  c = 32'he98fa333;
        7'b0110011 :  c = 32'he8dbf4fb;
        7'b0110100 :  c = 32'he82e0fa7;
        7'b0110101 :  c = 32'he7861eaf;
        7'b0110110 :  c = 32'he6e44c0f;
        7'b0110111 :  c = 32'he648c03a;
        7'b0111000 :  c = 32'he5b3a213;
        7'b0111001 :  c = 32'he52516e1;
        7'b0111010 :  c = 32'he49d4245;
        7'b0111011 :  c = 32'he41c4633;
        7'b0111100 :  c = 32'he3a242ec;
        7'b0111101 :  c = 32'he32f56ed;
        7'b0111110 :  c = 32'he2c39ef2;
        7'b0111111 :  c = 32'he25f35e9;
        7'b1000000 :  c = 32'he20234eb;
        7'b1000001 :  c = 32'he1acb337;
        7'b1000010 :  c = 32'he15ec62e;
        7'b1000011 :  c = 32'he118814b;
        7'b1000100 :  c = 32'he0d9f61e;
        7'b1000101 :  c = 32'he0a3344b;
        7'b1000110 :  c = 32'he0744980;
        7'b1000111 :  c = 32'he04d4179;
        7'b1001000 :  c = 32'he02e25f7;
        7'b1001001 :  c = 32'he016fec2;
        7'b1001010 :  c = 32'he007d1a2;
        7'b1001011 :  c = 32'he000a263;
        7'b1001100 :  c = 32'he00172d1;
        7'b1001101 :  c = 32'he00a42b7;
        7'b1001110 :  c = 32'he01b0fe2;
        7'b1001111 :  c = 32'he033d61f;
        7'b1010000 :  c = 32'he0548f3c;
        7'b1010001 :  c = 32'he07d330b;
        7'b1010010 :  c = 32'he0adb762;
        7'b1010011 :  c = 32'he0e61023;
        7'b1010100 :  c = 32'he1262f36;
        7'b1010101 :  c = 32'he16e0494;
        7'b1010110 :  c = 32'he1bd7e48;
        7'b1010111 :  c = 32'he2148874;
        7'b1011000 :  c = 32'he2730d56;
        7'b1011001 :  c = 32'he2d8f54d;
        7'b1011010 :  c = 32'he34626e0;
        7'b1011011 :  c = 32'he3ba86c3;
        7'b1011100 :  c = 32'he435f7df;
        7'b1011101 :  c = 32'he4b85b58;
        7'b1011110 :  c = 32'he5419095;
        7'b1011111 :  c = 32'he5d1754b;
        7'b1100000 :  c = 32'he667e581;
        7'b1100001 :  c = 32'he704bb9b;
        7'b1100010 :  c = 32'he7a7d065;
        7'b1100011 :  c = 32'he850fb1a;
        7'b1100100 :  c = 32'he9001171;
        7'b1100101 :  c = 32'he9b4e7a4;
        7'b1100110 :  c = 32'hea6f5081;
        7'b1100111 :  c = 32'heb2f1d6c;
        7'b1101000 :  c = 32'hebf41e74;
        7'b1101001 :  c = 32'hecbe225a;
        7'b1101010 :  c = 32'hed8cf69e;
        7'b1101011 :  c = 32'hee60678b;
        7'b1101100 :  c = 32'hef384047;
        7'b1101101 :  c = 32'hf0144add;
        7'b1101110 :  c = 32'hf0f4504a;
        7'b1101111 :  c = 32'hf1d81890;
        7'b1110000 :  c = 32'hf2bf6abc;
        7'b1110001 :  c = 32'hf3aa0cfc;
        7'b1110010 :  c = 32'hf497c4a9;
        7'b1110011 :  c = 32'hf5885655;
        7'b1110100 :  c = 32'hf67b85dd;
        7'b1110101 :  c = 32'hf7711678;
        7'b1110110 :  c = 32'hf868cac1;
        7'b1110111 :  c = 32'hf96264ce;
        7'b1111000 :  c = 32'hfa5da638;
        7'b1111001 :  c = 32'hfb5a5031;
        7'b1111010 :  c = 32'hfc582391;
        7'b1111011 :  c = 32'hfd56e0e2;
        7'b1111100 :  c = 32'hfe564878;
        7'b1111101 :  c = 32'hff561a79;
        7'b1111110 :  c = 32'h005616f3;
        7'b1111111 :  c = 32'h0155fde7;
        default    :  c = 'x;
    endcase

endmodule    
