`include "quadra.vh"

module lut
(
    input  x1_t  x1,
    output a_t   a,
    output b_t   b,
    output c_t   c
);
    // Read coefficients:
    always_comb
    unique casez (x1)
        7'b0000000 :  a = 25'h1a57d87;
        7'b0000001 :  a = 25'h1a85ccc;
        7'b0000010 :  a = 25'h1ab51fb;
        7'b0000011 :  a = 25'h1ae5c54;
        7'b0000100 :  a = 25'h1b17b15;
        7'b0000101 :  a = 25'h1b4ad78;
        7'b0000110 :  a = 25'h1b7f2ae;
        7'b0000111 :  a = 25'h1bb49e8;
        7'b0001000 :  a = 25'h1beb24e;
        7'b0001001 :  a = 25'h1c22b09;
        7'b0001010 :  a = 25'h1c5b337;
        7'b0001011 :  a = 25'h1c949f9;
        7'b0001100 :  a = 25'h1ccee68;
        7'b0001101 :  a = 25'h1d09f9b;
        7'b0001110 :  a = 25'h1d45ca6;
        7'b0001111 :  a = 25'h1d82499;
        7'b0010000 :  a = 25'h1dbf683;
        7'b0010001 :  a = 25'h1dfd170;
        7'b0010010 :  a = 25'h1e3b468;
        7'b0010011 :  a = 25'h1e79e72;
        7'b0010100 :  a = 25'h1eb8e95;
        7'b0010101 :  a = 25'h1ef83d4;
        7'b0010110 :  a = 25'h1f37d32;
        7'b0010111 :  a = 25'h1f779b1;
        7'b0011000 :  a = 25'h1fb7851;
        7'b0011001 :  a = 25'h1ff7813;
        7'b0011010 :  a = 25'h00377f6;
        7'b0011011 :  a = 25'h00776fc;
        7'b0011100 :  a = 25'h00b7425;
        7'b0011101 :  a = 25'h00f6e70;
        7'b0011110 :  a = 25'h01364e0;
        7'b0011111 :  a = 25'h0175677;
        7'b0100000 :  a = 25'h01b4238;
        7'b0100001 :  a = 25'h01f2729;
        7'b0100010 :  a = 25'h0230450;
        7'b0100011 :  a = 25'h026d8b6;
        7'b0100100 :  a = 25'h02aa367;
        7'b0100101 :  a = 25'h02e636e;
        7'b0100110 :  a = 25'h03217de;
        7'b0100111 :  a = 25'h035bfc7;
        7'b0101000 :  a = 25'h0395a41;
        7'b0101001 :  a = 25'h03ce664;
        7'b0101010 :  a = 25'h040634e;
        7'b0101011 :  a = 25'h043d020;
        7'b0101100 :  a = 25'h0472bfe;
        7'b0101101 :  a = 25'h04a7611;
        7'b0101110 :  a = 25'h04dad88;
        7'b0101111 :  a = 25'h050d193;
        7'b0110000 :  a = 25'h053e16b;
        7'b0110001 :  a = 25'h056dc4a;
        7'b0110010 :  a = 25'h059c173;
        7'b0110011 :  a = 25'h05c902b;
        7'b0110100 :  a = 25'h05f47c1;
        7'b0110101 :  a = 25'h061e785;
        7'b0110110 :  a = 25'h0646ecf;
        7'b0110111 :  a = 25'h066dcff;
        7'b0111000 :  a = 25'h0693177;
        7'b0111001 :  a = 25'h06b6ba4;
        7'b0111010 :  a = 25'h06d8af6;
        7'b0111011 :  a = 25'h06f8ee7;
        7'b0111100 :  a = 25'h07176f4;
        7'b0111101 :  a = 25'h07342a4;
        7'b0111110 :  a = 25'h074f184;
        7'b0111111 :  a = 25'h0768328;
        7'b1000000 :  a = 25'h077f72c;
        7'b1000001 :  a = 25'h0794d33;
        7'b1000010 :  a = 25'h07a84e7;
        7'b1000011 :  a = 25'h07b9dfa;
        7'b1000100 :  a = 25'h07c9827;
        7'b1000101 :  a = 25'h07d732e;
        7'b1000110 :  a = 25'h07e2ed9;
        7'b1000111 :  a = 25'h07ecafa;
        7'b1001000 :  a = 25'h07f4768;
        7'b1001001 :  a = 25'h07fa405;
        7'b1001010 :  a = 25'h07fe0b9;
        7'b1001011 :  a = 25'h07ffd76;
        7'b1001100 :  a = 25'h07ffa34;
        7'b1001101 :  a = 25'h07fd6f5;
        7'b1001110 :  a = 25'h07f93c0;
        7'b1001111 :  a = 25'h07f30a7;
        7'b1010000 :  a = 25'h07eadc3;
        7'b1010001 :  a = 25'h07e0b33;
        7'b1010010 :  a = 25'h07d4922;
        7'b1010011 :  a = 25'h07c67bf;
        7'b1010100 :  a = 25'h07b6743;
        7'b1010101 :  a = 25'h07a47ed;
        7'b1010110 :  a = 25'h0790a07;
        7'b1010111 :  a = 25'h077adde;
        7'b1011000 :  a = 25'h07633ca;
        7'b1011001 :  a = 25'h0749c2a;
        7'b1011010 :  a = 25'h072e764;
        7'b1011011 :  a = 25'h07115e5;
        7'b1011100 :  a = 25'h06f2820;
        7'b1011101 :  a = 25'h06d1e92;
        7'b1011110 :  a = 25'h06af9bd;
        7'b1011111 :  a = 25'h068ba2b;
        7'b1100000 :  a = 25'h066606a;
        7'b1100001 :  a = 25'h063ed11;
        7'b1100010 :  a = 25'h06160be;
        7'b1100011 :  a = 25'h05ebc13;
        7'b1100100 :  a = 25'h05bffba;
        7'b1100101 :  a = 25'h0592c61;
        7'b1100110 :  a = 25'h05642be;
        7'b1100111 :  a = 25'h053438a;
        7'b1101000 :  a = 25'h0502f86;
        7'b1101001 :  a = 25'h04d0777;
        7'b1101010 :  a = 25'h049cc25;
        7'b1101011 :  a = 25'h0467e62;
        7'b1101100 :  a = 25'h0431eff;
        7'b1101101 :  a = 25'h03faed4;
        7'b1101110 :  a = 25'h03c2ebf;
        7'b1101111 :  a = 25'h0389f9e;
        7'b1110000 :  a = 25'h0350255;
        7'b1110001 :  a = 25'h03157cc;
        7'b1110010 :  a = 25'h02da0ed;
        7'b1110011 :  a = 25'h029dea7;
        7'b1110100 :  a = 25'h02611e8;
        7'b1110101 :  a = 25'h0223ba6;
        7'b1110110 :  a = 25'h01e5cd5;
        7'b1110111 :  a = 25'h01a766d;
        7'b1111000 :  a = 25'h0168967;
        7'b1111001 :  a = 25'h01296bf;
        7'b1111010 :  a = 25'h00e9f72;
        7'b1111011 :  a = 25'h00aa47c;
        7'b1111100 :  a = 25'h006a6de;
        7'b1111101 :  a = 25'h002a796;
        7'b1111110 :  a = 25'h1fea7a5;
        7'b1111111 :  a = 25'h1faa809;
        default    :  a = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  b = 19'h16a0c;
        7'b0000001 :  b = 19'h1752f;
        7'b0000010 :  b = 19'h17ff4;
        7'b0000011 :  b = 19'h18a59;
        7'b0000100 :  b = 19'h1945c;
        7'b0000101 :  b = 19'h19dfa;
        7'b0000110 :  b = 19'h1a730;
        7'b0000111 :  b = 19'h1affd;
        7'b0001000 :  b = 19'h1b85d;
        7'b0001001 :  b = 19'h1c04f;
        7'b0001010 :  b = 19'h1c7d2;
        7'b0001011 :  b = 19'h1cee2;
        7'b0001100 :  b = 19'h1d57f;
        7'b0001101 :  b = 19'h1dba6;
        7'b0001110 :  b = 19'h1e156;
        7'b0001111 :  b = 19'h1e68e;
        7'b0010000 :  b = 19'h1eb4d;
        7'b0010001 :  b = 19'h1ef91;
        7'b0010010 :  b = 19'h1f358;
        7'b0010011 :  b = 19'h1f6a3;
        7'b0010100 :  b = 19'h1f970;
        7'b0010101 :  b = 19'h1fbbf;
        7'b0010110 :  b = 19'h1fd8f;
        7'b0010111 :  b = 19'h1fee0;
        7'b0011000 :  b = 19'h1ffb1;
        7'b0011001 :  b = 19'h20002;
        7'b0011010 :  b = 19'h1ffd3;
        7'b0011011 :  b = 19'h1ff24;
        7'b0011100 :  b = 19'h1fdf5;
        7'b0011101 :  b = 19'h1fc47;
        7'b0011110 :  b = 19'h1fa1a;
        7'b0011111 :  b = 19'h1f76e;
        7'b0100000 :  b = 19'h1f444;
        7'b0100001 :  b = 19'h1f09e;
        7'b0100010 :  b = 19'h1ec7b;
        7'b0100011 :  b = 19'h1e7dd;
        7'b0100100 :  b = 19'h1e2c5;
        7'b0100101 :  b = 19'h1dd34;
        7'b0100110 :  b = 19'h1d72c;
        7'b0100111 :  b = 19'h1d0af;
        7'b0101000 :  b = 19'h1c9bd;
        7'b0101001 :  b = 19'h1c259;
        7'b0101010 :  b = 19'h1ba84;
        7'b0101011 :  b = 19'h1b240;
        7'b0101100 :  b = 19'h1a990;
        7'b0101101 :  b = 19'h1a076;
        7'b0101110 :  b = 19'h196f4;
        7'b0101111 :  b = 19'h18d0b;
        7'b0110000 :  b = 19'h182c0;
        7'b0110001 :  b = 19'h17814;
        7'b0110010 :  b = 19'h16d0a;
        7'b0110011 :  b = 19'h161a4;
        7'b0110100 :  b = 19'h155e6;
        7'b0110101 :  b = 19'h149d3;
        7'b0110110 :  b = 19'h13d6d;
        7'b0110111 :  b = 19'h130b8;
        7'b0111000 :  b = 19'h123b7;
        7'b0111001 :  b = 19'h1166d;
        7'b0111010 :  b = 19'h108dd;
        7'b0111011 :  b = 19'h0fb0b;
        7'b0111100 :  b = 19'h0ecfa;
        7'b0111101 :  b = 19'h0deae;
        7'b0111110 :  b = 19'h0d02b;
        7'b0111111 :  b = 19'h0c173;
        7'b1000000 :  b = 19'h0b28b;
        7'b1000001 :  b = 19'h0a376;
        7'b1000010 :  b = 19'h09439;
        7'b1000011 :  b = 19'h084d6;
        7'b1000100 :  b = 19'h07552;
        7'b1000101 :  b = 19'h065b1;
        7'b1000110 :  b = 19'h055f7;
        7'b1000111 :  b = 19'h04627;
        7'b1001000 :  b = 19'h03645;
        7'b1001001 :  b = 19'h02656;
        7'b1001010 :  b = 19'h0165d;
        7'b1001011 :  b = 19'h0065f;
        7'b1001100 :  b = 19'h7f65f;
        7'b1001101 :  b = 19'h7e662;
        7'b1001110 :  b = 19'h7d66b;
        7'b1001111 :  b = 19'h7c67e;
        7'b1010000 :  b = 19'h7b6a0;
        7'b1010001 :  b = 19'h7a6d4;
        7'b1010010 :  b = 19'h7971e;
        7'b1010011 :  b = 19'h78783;
        7'b1010100 :  b = 19'h77805;
        7'b1010101 :  b = 19'h768aa;
        7'b1010110 :  b = 19'h75974;
        7'b1010111 :  b = 19'h74a68;
        7'b1011000 :  b = 19'h73b8a;
        7'b1011001 :  b = 19'h72cdd;
        7'b1011010 :  b = 19'h71e64;
        7'b1011011 :  b = 19'h71024;
        7'b1011100 :  b = 19'h7021f;
        7'b1011101 :  b = 19'h6f45b;
        7'b1011110 :  b = 19'h6e6d9;
        7'b1011111 :  b = 19'h6d99d;
        7'b1100000 :  b = 19'h6ccab;
        7'b1100001 :  b = 19'h6c006;
        7'b1100010 :  b = 19'h6b3b1;
        7'b1100011 :  b = 19'h6a7af;
        7'b1100100 :  b = 19'h69c03;
        7'b1100101 :  b = 19'h690b0;
        7'b1100110 :  b = 19'h685b8;
        7'b1100111 :  b = 19'h67b20;
        7'b1101000 :  b = 19'h670e8;
        7'b1101001 :  b = 19'h66714;
        7'b1101010 :  b = 19'h65da7;
        7'b1101011 :  b = 19'h654a2;
        7'b1101100 :  b = 19'h64c08;
        7'b1101101 :  b = 19'h643db;
        7'b1101110 :  b = 19'h63c1d;
        7'b1101111 :  b = 19'h634d0;
        7'b1110000 :  b = 19'h62df5;
        7'b1110001 :  b = 19'h62790;
        7'b1110010 :  b = 19'h621a0;
        7'b1110011 :  b = 19'h61c28;
        7'b1110100 :  b = 19'h61729;
        7'b1110101 :  b = 19'h612a4;
        7'b1110110 :  b = 19'h60e9a;
        7'b1110111 :  b = 19'h60b0d;
        7'b1111000 :  b = 19'h607fd;
        7'b1111001 :  b = 19'h6056b;
        7'b1111010 :  b = 19'h60357;
        7'b1111011 :  b = 19'h601c3;
        7'b1111100 :  b = 19'h600ae;
        7'b1111101 :  b = 19'h60019;
        7'b1111110 :  b = 19'h60004;
        7'b1111111 :  b = 19'h6006f;
        default    :  b = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  c = 15'h2ce6;
        7'b0000001 :  c = 15'h2b74;
        7'b0000010 :  c = 15'h29f6;
        7'b0000011 :  c = 15'h286e;
        7'b0000100 :  c = 15'h26de;
        7'b0000101 :  c = 15'h2542;
        7'b0000110 :  c = 15'h239c;
        7'b0000111 :  c = 15'h21ee;
        7'b0001000 :  c = 15'h2038;
        7'b0001001 :  c = 15'h1e7a;
        7'b0001010 :  c = 15'h1cb4;
        7'b0001011 :  c = 15'h1ae8;
        7'b0001100 :  c = 15'h1914;
        7'b0001101 :  c = 15'h173a;
        7'b0001110 :  c = 15'h155a;
        7'b0001111 :  c = 15'h1374;
        7'b0010000 :  c = 15'h118a;
        7'b0010001 :  c = 15'h0f9c;
        7'b0010010 :  c = 15'h0da8;
        7'b0010011 :  c = 15'h0bb4;
        7'b0010100 :  c = 15'h09ba;
        7'b0010101 :  c = 15'h07c0;
        7'b0010110 :  c = 15'h05c2;
        7'b0010111 :  c = 15'h03c4;
        7'b0011000 :  c = 15'h01c4;
        7'b0011001 :  c = 15'h7fc4;
        7'b0011010 :  c = 15'h7dc4;
        7'b0011011 :  c = 15'h7bc4;
        7'b0011100 :  c = 15'h79c6;
        7'b0011101 :  c = 15'h77ca;
        7'b0011110 :  c = 15'h75d0;
        7'b0011111 :  c = 15'h73d8;
        7'b0100000 :  c = 15'h71e2;
        7'b0100001 :  c = 15'h6ff0;
        7'b0100010 :  c = 15'h6e02;
        7'b0100011 :  c = 15'h6c1a;
        7'b0100100 :  c = 15'h6a36;
        7'b0100101 :  c = 15'h6858;
        7'b0100110 :  c = 15'h667e;
        7'b0100111 :  c = 15'h64ac;
        7'b0101000 :  c = 15'h62e0;
        7'b0101001 :  c = 15'h611c;
        7'b0101010 :  c = 15'h5f60;
        7'b0101011 :  c = 15'h5dac;
        7'b0101100 :  c = 15'h5c00;
        7'b0101101 :  c = 15'h5a5e;
        7'b0101110 :  c = 15'h58c4;
        7'b0101111 :  c = 15'h5734;
        7'b0110000 :  c = 15'h55ae;
        7'b0110001 :  c = 15'h5434;
        7'b0110010 :  c = 15'h52c4;
        7'b0110011 :  c = 15'h5160;
        7'b0110100 :  c = 15'h5008;
        7'b0110101 :  c = 15'h4eba;
        7'b0110110 :  c = 15'h4d7a;
        7'b0110111 :  c = 15'h4c46;
        7'b0111000 :  c = 15'h4b1e;
        7'b0111001 :  c = 15'h4a06;
        7'b0111010 :  c = 15'h48f8;
        7'b0111011 :  c = 15'h47fa;
        7'b0111100 :  c = 15'h470a;
        7'b0111101 :  c = 15'h4628;
        7'b0111110 :  c = 15'h4554;
        7'b0111111 :  c = 15'h448e;
        7'b1000000 :  c = 15'h43d8;
        7'b1000001 :  c = 15'h4332;
        7'b1000010 :  c = 15'h429a;
        7'b1000011 :  c = 15'h4210;
        7'b1000100 :  c = 15'h4198;
        7'b1000101 :  c = 15'h412e;
        7'b1000110 :  c = 15'h40d4;
        7'b1000111 :  c = 15'h408a;
        7'b1001000 :  c = 15'h4050;
        7'b1001001 :  c = 15'h4024;
        7'b1001010 :  c = 15'h400a;
        7'b1001011 :  c = 15'h4000;
        7'b1001100 :  c = 15'h4006;
        7'b1001101 :  c = 15'h401c;
        7'b1001110 :  c = 15'h4042;
        7'b1001111 :  c = 15'h4076;
        7'b1010000 :  c = 15'h40bc;
        7'b1010001 :  c = 15'h4112;
        7'b1010010 :  c = 15'h4176;
        7'b1010011 :  c = 15'h41ea;
        7'b1010100 :  c = 15'h426e;
        7'b1010101 :  c = 15'h4302;
        7'b1010110 :  c = 15'h43a6;
        7'b1010111 :  c = 15'h4456;
        7'b1011000 :  c = 15'h4518;
        7'b1011001 :  c = 15'h45e8;
        7'b1011010 :  c = 15'h46c6;
        7'b1011011 :  c = 15'h47b2;
        7'b1011100 :  c = 15'h48ac;
        7'b1011101 :  c = 15'h49b4;
        7'b1011110 :  c = 15'h4aca;
        7'b1011111 :  c = 15'h4bec;
        7'b1100000 :  c = 15'h4d1e;
        7'b1100001 :  c = 15'h4e5a;
        7'b1100010 :  c = 15'h4fa4;
        7'b1100011 :  c = 15'h50f8;
        7'b1100100 :  c = 15'h525a;
        7'b1100101 :  c = 15'h53c6;
        7'b1100110 :  c = 15'h553e;
        7'b1100111 :  c = 15'h56c0;
        7'b1101000 :  c = 15'h584c;
        7'b1101001 :  c = 15'h59e2;
        7'b1101010 :  c = 15'h5b82;
        7'b1101011 :  c = 15'h5d2c;
        7'b1101100 :  c = 15'h5ede;
        7'b1101101 :  c = 15'h6098;
        7'b1101110 :  c = 15'h625a;
        7'b1101111 :  c = 15'h6424;
        7'b1110000 :  c = 15'h65f4;
        7'b1110001 :  c = 15'h67ca;
        7'b1110010 :  c = 15'h69a8;
        7'b1110011 :  c = 15'h6b8a;
        7'b1110100 :  c = 15'h6d72;
        7'b1110101 :  c = 15'h6f5e;
        7'b1110110 :  c = 15'h714e;
        7'b1110111 :  c = 15'h7342;
        7'b1111000 :  c = 15'h753a;
        7'b1111001 :  c = 15'h7734;
        7'b1111010 :  c = 15'h7930;
        7'b1111011 :  c = 15'h7b2e;
        7'b1111100 :  c = 15'h7d2c;
        7'b1111101 :  c = 15'h7f2c;
        7'b1111110 :  c = 15'h012c;
        7'b1111111 :  c = 15'h032c;
        default    :  c = 'x;
    endcase

endmodule
