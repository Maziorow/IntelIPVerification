`include "quadra.vh"

module lut
(
    input  x1_t  x1,
    output a_t   a,
    output b_t   b,
    output c_t   c
);
    // Read coefficients:
    always_comb
    unique casez (x1)
        7'b0000000 :  a = 27'h695f619;
        7'b0000001 :  a = 27'h6a17330;
        7'b0000010 :  a = 27'h6ad47e9;
        7'b0000011 :  a = 27'h6b9714d;
        7'b0000100 :  a = 27'h6c5ec53;
        7'b0000101 :  a = 27'h6d2b5dd;
        7'b0000110 :  a = 27'h6dfcab7;
        7'b0000111 :  a = 27'h6ed279d;
        7'b0001000 :  a = 27'h6fac938;
        7'b0001001 :  a = 27'h708ac21;
        7'b0001010 :  a = 27'h716ccdb;
        7'b0001011 :  a = 27'h72527e2;
        7'b0001100 :  a = 27'h733b99e;
        7'b0001101 :  a = 27'h7427e6a;
        7'b0001110 :  a = 27'h7517296;
        7'b0001111 :  a = 27'h7609264;
        7'b0010000 :  a = 27'h76fda0c;
        7'b0010001 :  a = 27'h77f45bd;
        7'b0010010 :  a = 27'h78ed19d;
        7'b0010011 :  a = 27'h79e79c7;
        7'b0010100 :  a = 27'h7ae3a53;
        7'b0010101 :  a = 27'h7be0f4f;
        7'b0010110 :  a = 27'h7cdf4c7;
        7'b0010111 :  a = 27'h7dde6c2;
        7'b0011000 :  a = 27'h7ede142;
        7'b0011001 :  a = 27'h7fde04a;
        7'b0011010 :  a = 27'h00ddfda;
        7'b0011011 :  a = 27'h01ddbf3;
        7'b0011100 :  a = 27'h02dd094;
        7'b0011101 :  a = 27'h03db9c2;
        7'b0011110 :  a = 27'h04d9381;
        7'b0011111 :  a = 27'h05d59dc;
        7'b0100000 :  a = 27'h06d08e1;
        7'b0100001 :  a = 27'h07c9ca4;
        7'b0100010 :  a = 27'h08c1142;
        7'b0100011 :  a = 27'h09b62db;
        7'b0100100 :  a = 27'h0aa8d9d;
        7'b0100101 :  a = 27'h0b98dbb;
        7'b0100110 :  a = 27'h0c85f78;
        7'b0100111 :  a = 27'h0d6ff1e;
        7'b0101000 :  a = 27'h0e56905;
        7'b0101001 :  a = 27'h0f39992;
        7'b0101010 :  a = 27'h1018d3b;
        7'b0101011 :  a = 27'h10f4082;
        7'b0101100 :  a = 27'h11caffa;
        7'b0101101 :  a = 27'h129d847;
        7'b0101110 :  a = 27'h136b620;
        7'b0101111 :  a = 27'h143464e;
        7'b0110000 :  a = 27'h14f85ac;
        7'b0110001 :  a = 27'h15b7129;
        7'b0110010 :  a = 27'h16705cc;
        7'b0110011 :  a = 27'h17240af;
        7'b0110100 :  a = 27'h17d1f05;
        7'b0110101 :  a = 27'h1879e14;
        7'b0110110 :  a = 27'h191bb3e;
        7'b0110111 :  a = 27'h19b73fc;
        7'b0111000 :  a = 27'h1a4c5de;
        7'b0111001 :  a = 27'h1adae91;
        7'b0111010 :  a = 27'h1b62bdb;
        7'b0111011 :  a = 27'h1be3b9c;
        7'b0111100 :  a = 27'h1c5dbd1;
        7'b0111101 :  a = 27'h1cd0a91;
        7'b0111110 :  a = 27'h1d3c610;
        7'b0111111 :  a = 27'h1da0ca0;
        7'b1000000 :  a = 27'h1dfdcb1;
        7'b1000001 :  a = 27'h1e534cc;
        7'b1000010 :  a = 27'h1ea139c;
        7'b1000011 :  a = 27'h1ee77eb;
        7'b1000100 :  a = 27'h1f2609e;
        7'b1000101 :  a = 27'h1f5ccbb;
        7'b1000110 :  a = 27'h1f8bb67;
        7'b1000111 :  a = 27'h1fb2be8;
        7'b1001000 :  a = 27'h1fd1da0;
        7'b1001001 :  a = 27'h1fe9014;
        7'b1001010 :  a = 27'h1ff82e6;
        7'b1001011 :  a = 27'h1fff5da;
        7'b1001100 :  a = 27'h1ffe8d3;
        7'b1001101 :  a = 27'h1ff5bd5;
        7'b1001110 :  a = 27'h1fe4f02;
        7'b1001111 :  a = 27'h1fcc29e;
        7'b1010000 :  a = 27'h1fab70c;
        7'b1010001 :  a = 27'h1f82ccf;
        7'b1010010 :  a = 27'h1f5248a;
        7'b1010011 :  a = 27'h1f19efe;
        7'b1010100 :  a = 27'h1ed9d0d;
        7'b1010101 :  a = 27'h1e91fb7;
        7'b1010110 :  a = 27'h1e4281c;
        7'b1010111 :  a = 27'h1deb779;
        7'b1011000 :  a = 27'h1d8cf2b;
        7'b1011001 :  a = 27'h1d270ab;
        7'b1011010 :  a = 27'h1cb9d93;
        7'b1011011 :  a = 27'h1c45794;
        7'b1011100 :  a = 27'h1bca083;
        7'b1011101 :  a = 27'h1b47a4b;
        7'b1011110 :  a = 27'h1abe6f7;
        7'b1011111 :  a = 27'h1a2e8ac;
        7'b1100000 :  a = 27'h19981a8;
        7'b1100001 :  a = 27'h18fb446;
        7'b1100010 :  a = 27'h18582fa;
        7'b1100011 :  a = 27'h17af04f;
        7'b1100100 :  a = 27'h16ffee9;
        7'b1100101 :  a = 27'h164b186;
        7'b1100110 :  a = 27'h1590af9;
        7'b1100111 :  a = 27'h14d0e2a;
        7'b1101000 :  a = 27'h140be19;
        7'b1101001 :  a = 27'h1341ddc;
        7'b1101010 :  a = 27'h1273096;
        7'b1101011 :  a = 27'h119f988;
        7'b1101100 :  a = 27'h10c7bfc;
        7'b1101101 :  a = 27'h0febb53;
        7'b1101110 :  a = 27'h0f0bafc;
        7'b1101111 :  a = 27'h0e27e78;
        7'b1110000 :  a = 27'h0d40955;
        7'b1110001 :  a = 27'h0c55f31;
        7'b1110010 :  a = 27'h0b683b7;
        7'b1110011 :  a = 27'h0a77a9c;
        7'b1110100 :  a = 27'h09847a3;
        7'b1110101 :  a = 27'h088ee99;
        7'b1110110 :  a = 27'h0797354;
        7'b1110111 :  a = 27'h069d9b4;
        7'b1111000 :  a = 27'h05a259d;
        7'b1111001 :  a = 27'h04a5afd;
        7'b1111010 :  a = 27'h03a7dc8;
        7'b1111011 :  a = 27'h02a91f3;
        7'b1111100 :  a = 27'h01a9b79;
        7'b1111101 :  a = 27'h00a9e59;
        7'b1111110 :  a = 27'h7fa9e92;
        7'b1111111 :  a = 27'h7eaa023;
        default    :  a = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  b = 20'h2d418;
        7'b0000001 :  b = 20'h2ea5e;
        7'b0000010 :  b = 20'h2ffe8;
        7'b0000011 :  b = 20'h314b3;
        7'b0000100 :  b = 20'h328b9;
        7'b0000101 :  b = 20'h33bf4;
        7'b0000110 :  b = 20'h34e61;
        7'b0000111 :  b = 20'h35ffa;
        7'b0001000 :  b = 20'h370bb;
        7'b0001001 :  b = 20'h3809f;
        7'b0001010 :  b = 20'h38fa4;
        7'b0001011 :  b = 20'h39dc5;
        7'b0001100 :  b = 20'h3aafe;
        7'b0001101 :  b = 20'h3b74d;
        7'b0001110 :  b = 20'h3c2ad;
        7'b0001111 :  b = 20'h3cd1d;
        7'b0010000 :  b = 20'h3d69a;
        7'b0010001 :  b = 20'h3df22;
        7'b0010010 :  b = 20'h3e6b1;
        7'b0010011 :  b = 20'h3ed47;
        7'b0010100 :  b = 20'h3f2e1;
        7'b0010101 :  b = 20'h3f77f;
        7'b0010110 :  b = 20'h3fb1f;
        7'b0010111 :  b = 20'h3fdc0;
        7'b0011000 :  b = 20'h3ff62;
        7'b0011001 :  b = 20'h40004;
        7'b0011010 :  b = 20'h3ffa6;
        7'b0011011 :  b = 20'h3fe48;
        7'b0011100 :  b = 20'h3fbeb;
        7'b0011101 :  b = 20'h3f88e;
        7'b0011110 :  b = 20'h3f434;
        7'b0011111 :  b = 20'h3eedc;
        7'b0100000 :  b = 20'h3e889;
        7'b0100001 :  b = 20'h3e13c;
        7'b0100010 :  b = 20'h3d8f6;
        7'b0100011 :  b = 20'h3cfba;
        7'b0100100 :  b = 20'h3c58a;
        7'b0100101 :  b = 20'h3ba69;
        7'b0100110 :  b = 20'h3ae59;
        7'b0100111 :  b = 20'h3a15e;
        7'b0101000 :  b = 20'h3937a;
        7'b0101001 :  b = 20'h384b2;
        7'b0101010 :  b = 20'h37508;
        7'b0101011 :  b = 20'h36481;
        7'b0101100 :  b = 20'h35321;
        7'b0101101 :  b = 20'h340ed;
        7'b0101110 :  b = 20'h32de8;
        7'b0101111 :  b = 20'h31a17;
        7'b0110000 :  b = 20'h30580;
        7'b0110001 :  b = 20'h2f028;
        7'b0110010 :  b = 20'h2da14;
        7'b0110011 :  b = 20'h2c349;
        7'b0110100 :  b = 20'h2abcd;
        7'b0110101 :  b = 20'h293a7;
        7'b0110110 :  b = 20'h27adb;
        7'b0110111 :  b = 20'h26171;
        7'b0111000 :  b = 20'h2476f;
        7'b0111001 :  b = 20'h22cda;
        7'b0111010 :  b = 20'h211bb;
        7'b0111011 :  b = 20'h1f617;
        7'b0111100 :  b = 20'h1d9f5;
        7'b0111101 :  b = 20'h1bd5d;
        7'b0111110 :  b = 20'h1a056;
        7'b0111111 :  b = 20'h182e7;
        7'b1000000 :  b = 20'h16516;
        7'b1000001 :  b = 20'h146ed;
        7'b1000010 :  b = 20'h12872;
        7'b1000011 :  b = 20'h109ad;
        7'b1000100 :  b = 20'h0eaa5;
        7'b1000101 :  b = 20'h0cb63;
        7'b1000110 :  b = 20'h0abee;
        7'b1000111 :  b = 20'h08c4e;
        7'b1001000 :  b = 20'h06c8b;
        7'b1001001 :  b = 20'h04cac;
        7'b1001010 :  b = 20'h02cbb;
        7'b1001011 :  b = 20'h00cbe;
        7'b1001100 :  b = 20'hfecbe;
        7'b1001101 :  b = 20'hfccc3;
        7'b1001110 :  b = 20'hfacd5;
        7'b1001111 :  b = 20'hf8cfc;
        7'b1010000 :  b = 20'hf6d3f;
        7'b1010001 :  b = 20'hf4da7;
        7'b1010010 :  b = 20'hf2e3c;
        7'b1010011 :  b = 20'hf0f05;
        7'b1010100 :  b = 20'hef00a;
        7'b1010101 :  b = 20'hed153;
        7'b1010110 :  b = 20'heb2e8;
        7'b1010111 :  b = 20'he94d0;
        7'b1011000 :  b = 20'he7713;
        7'b1011001 :  b = 20'he59b9;
        7'b1011010 :  b = 20'he3cc7;
        7'b1011011 :  b = 20'he2047;
        7'b1011100 :  b = 20'he043e;
        7'b1011101 :  b = 20'hde8b5;
        7'b1011110 :  b = 20'hdcdb1;
        7'b1011111 :  b = 20'hdb33a;
        7'b1100000 :  b = 20'hd9956;
        7'b1100001 :  b = 20'hd800c;
        7'b1100010 :  b = 20'hd6761;
        7'b1100011 :  b = 20'hd4f5d;
        7'b1100100 :  b = 20'hd3805;
        7'b1100101 :  b = 20'hd215f;
        7'b1100110 :  b = 20'hd0b70;
        7'b1100111 :  b = 20'hcf63f;
        7'b1101000 :  b = 20'hce1d0;
        7'b1101001 :  b = 20'hcce28;
        7'b1101010 :  b = 20'hcbb4e;
        7'b1101011 :  b = 20'hca944;
        7'b1101100 :  b = 20'hc9810;
        7'b1101101 :  b = 20'hc87b5;
        7'b1101110 :  b = 20'hc7839;
        7'b1101111 :  b = 20'hc699f;
        7'b1110000 :  b = 20'hc5bea;
        7'b1110001 :  b = 20'hc4f1f;
        7'b1110010 :  b = 20'hc433f;
        7'b1110011 :  b = 20'hc384f;
        7'b1110100 :  b = 20'hc2e51;
        7'b1110101 :  b = 20'hc2547;
        7'b1110110 :  b = 20'hc1d34;
        7'b1110111 :  b = 20'hc1619;
        7'b1111000 :  b = 20'hc0ff9;
        7'b1111001 :  b = 20'hc0ad5;
        7'b1111010 :  b = 20'hc06ae;
        7'b1111011 :  b = 20'hc0385;
        7'b1111100 :  b = 20'hc015c;
        7'b1111101 :  b = 20'hc0032;
        7'b1111110 :  b = 20'hc0008;
        7'b1111111 :  b = 20'hc00de;
        default    :  b = 'x;
    endcase

    always_comb
    unique casez (x1)
        7'b0000000 :  c = 16'h59cc;
        7'b0000001 :  c = 16'h56e8;
        7'b0000010 :  c = 16'h53ec;
        7'b0000011 :  c = 16'h50dc;
        7'b0000100 :  c = 16'h4dbc;
        7'b0000101 :  c = 16'h4a84;
        7'b0000110 :  c = 16'h4738;
        7'b0000111 :  c = 16'h43dc;
        7'b0001000 :  c = 16'h4070;
        7'b0001001 :  c = 16'h3cf4;
        7'b0001010 :  c = 16'h3968;
        7'b0001011 :  c = 16'h35d0;
        7'b0001100 :  c = 16'h3228;
        7'b0001101 :  c = 16'h2e74;
        7'b0001110 :  c = 16'h2ab4;
        7'b0001111 :  c = 16'h26e8;
        7'b0010000 :  c = 16'h2314;
        7'b0010001 :  c = 16'h1f38;
        7'b0010010 :  c = 16'h1b50;
        7'b0010011 :  c = 16'h1768;
        7'b0010100 :  c = 16'h1374;
        7'b0010101 :  c = 16'h0f80;
        7'b0010110 :  c = 16'h0b84;
        7'b0010111 :  c = 16'h0788;
        7'b0011000 :  c = 16'h0388;
        7'b0011001 :  c = 16'hff88;
        7'b0011010 :  c = 16'hfb88;
        7'b0011011 :  c = 16'hf788;
        7'b0011100 :  c = 16'hf38c;
        7'b0011101 :  c = 16'hef94;
        7'b0011110 :  c = 16'heba0;
        7'b0011111 :  c = 16'he7b0;
        7'b0100000 :  c = 16'he3c4;
        7'b0100001 :  c = 16'hdfe0;
        7'b0100010 :  c = 16'hdc04;
        7'b0100011 :  c = 16'hd834;
        7'b0100100 :  c = 16'hd46c;
        7'b0100101 :  c = 16'hd0b0;
        7'b0100110 :  c = 16'hccfc;
        7'b0100111 :  c = 16'hc958;
        7'b0101000 :  c = 16'hc5c0;
        7'b0101001 :  c = 16'hc238;
        7'b0101010 :  c = 16'hbec0;
        7'b0101011 :  c = 16'hbb58;
        7'b0101100 :  c = 16'hb800;
        7'b0101101 :  c = 16'hb4bc;
        7'b0101110 :  c = 16'hb188;
        7'b0101111 :  c = 16'hae68;
        7'b0110000 :  c = 16'hab5c;
        7'b0110001 :  c = 16'ha868;
        7'b0110010 :  c = 16'ha588;
        7'b0110011 :  c = 16'ha2c0;
        7'b0110100 :  c = 16'ha010;
        7'b0110101 :  c = 16'h9d74;
        7'b0110110 :  c = 16'h9af4;
        7'b0110111 :  c = 16'h988c;
        7'b0111000 :  c = 16'h963c;
        7'b0111001 :  c = 16'h940c;
        7'b0111010 :  c = 16'h91f0;
        7'b0111011 :  c = 16'h8ff4;
        7'b0111100 :  c = 16'h8e14;
        7'b0111101 :  c = 16'h8c50;
        7'b0111110 :  c = 16'h8aa8;
        7'b0111111 :  c = 16'h891c;
        7'b1000000 :  c = 16'h87b0;
        7'b1000001 :  c = 16'h8664;
        7'b1000010 :  c = 16'h8534;
        7'b1000011 :  c = 16'h8420;
        7'b1000100 :  c = 16'h8330;
        7'b1000101 :  c = 16'h825c;
        7'b1000110 :  c = 16'h81a8;
        7'b1000111 :  c = 16'h8114;
        7'b1001000 :  c = 16'h80a0;
        7'b1001001 :  c = 16'h8048;
        7'b1001010 :  c = 16'h8014;
        7'b1001011 :  c = 16'h8000;
        7'b1001100 :  c = 16'h800c;
        7'b1001101 :  c = 16'h8038;
        7'b1001110 :  c = 16'h8084;
        7'b1001111 :  c = 16'h80ec;
        7'b1010000 :  c = 16'h8178;
        7'b1010001 :  c = 16'h8224;
        7'b1010010 :  c = 16'h82ec;
        7'b1010011 :  c = 16'h83d4;
        7'b1010100 :  c = 16'h84dc;
        7'b1010101 :  c = 16'h8604;
        7'b1010110 :  c = 16'h874c;
        7'b1010111 :  c = 16'h88ac;
        7'b1011000 :  c = 16'h8a30;
        7'b1011001 :  c = 16'h8bd0;
        7'b1011010 :  c = 16'h8d8c;
        7'b1011011 :  c = 16'h8f64;
        7'b1011100 :  c = 16'h9158;
        7'b1011101 :  c = 16'h9368;
        7'b1011110 :  c = 16'h9594;
        7'b1011111 :  c = 16'h97d8;
        7'b1100000 :  c = 16'h9a3c;
        7'b1100001 :  c = 16'h9cb4;
        7'b1100010 :  c = 16'h9f48;
        7'b1100011 :  c = 16'ha1f0;
        7'b1100100 :  c = 16'ha4b4;
        7'b1100101 :  c = 16'ha78c;
        7'b1100110 :  c = 16'haa7c;
        7'b1100111 :  c = 16'had80;
        7'b1101000 :  c = 16'hb098;
        7'b1101001 :  c = 16'hb3c4;
        7'b1101010 :  c = 16'hb704;
        7'b1101011 :  c = 16'hba58;
        7'b1101100 :  c = 16'hbdbc;
        7'b1101101 :  c = 16'hc130;
        7'b1101110 :  c = 16'hc4b4;
        7'b1101111 :  c = 16'hc848;
        7'b1110000 :  c = 16'hcbe8;
        7'b1110001 :  c = 16'hcf94;
        7'b1110010 :  c = 16'hd350;
        7'b1110011 :  c = 16'hd714;
        7'b1110100 :  c = 16'hdae4;
        7'b1110101 :  c = 16'hdebc;
        7'b1110110 :  c = 16'he29c;
        7'b1110111 :  c = 16'he684;
        7'b1111000 :  c = 16'hea74;
        7'b1111001 :  c = 16'hee68;
        7'b1111010 :  c = 16'hf260;
        7'b1111011 :  c = 16'hf65c;
        7'b1111100 :  c = 16'hfa58;
        7'b1111101 :  c = 16'hfe58;
        7'b1111110 :  c = 16'h0258;
        7'b1111111 :  c = 16'h0658;
        default    :  c = 'x;
    endcase

endmodule
